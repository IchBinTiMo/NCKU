module Decoder (
  ports
);
  
endmodule